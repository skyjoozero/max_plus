library verilog;
use verilog.vl_types.all;
entity example_vlg_vec_tst is
end example_vlg_vec_tst;
