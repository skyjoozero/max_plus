library verilog;
use verilog.vl_types.all;
entity dff_single_vlg_vec_tst is
end dff_single_vlg_vec_tst;
