library verilog;
use verilog.vl_types.all;
entity test is
    port(
        and2_out        : out    vl_logic;
        in0             : in     vl_logic;
        in1             : in     vl_logic
    );
end test;
