library verilog;
use verilog.vl_types.all;
entity dff_double_vlg_vec_tst is
end dff_double_vlg_vec_tst;
